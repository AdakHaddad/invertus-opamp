magic
tech sky130A
magscale 1 2
timestamp 1729350307
<< nwell >>
rect -206 -342 672 2046
<< nsubdiff >>
rect -170 1976 -110 2010
rect 576 1976 636 2010
rect -170 1945 -136 1976
rect 602 1945 636 1976
rect -170 -269 -136 -243
rect 602 -269 636 -243
rect -170 -303 -110 -269
rect 576 -303 636 -269
<< nsubdiffcont >>
rect -110 1976 576 2010
rect -170 -243 -136 1945
rect 602 -243 636 1945
rect -110 -303 576 -269
<< poly >>
rect 6 1448 36 1479
rect -54 1432 36 1448
rect -54 1398 -38 1432
rect -4 1398 36 1432
rect 410 1448 440 1489
rect 410 1432 500 1448
rect 410 1398 450 1432
rect 484 1398 500 1432
rect -54 1382 12 1398
rect 434 1382 500 1398
rect 6 954 36 984
rect -54 938 36 954
rect -54 904 -38 938
rect -4 904 36 938
rect 410 954 440 985
rect 410 938 500 954
rect 410 904 450 938
rect 484 904 500 938
rect -54 888 12 904
rect 434 888 500 904
rect 94 788 194 888
rect 252 788 352 888
rect -54 772 12 788
rect 434 772 500 788
rect -54 738 -38 772
rect -4 738 36 772
rect -54 722 36 738
rect 6 691 36 722
rect 410 738 450 772
rect 484 738 500 772
rect 410 722 500 738
rect 410 692 440 722
rect -54 278 12 294
rect 434 278 500 294
rect -54 244 -38 278
rect -4 244 36 278
rect -54 228 36 244
rect 6 197 36 228
rect 410 244 450 278
rect 484 244 500 278
rect 410 228 500 244
rect 410 198 440 228
<< polycont >>
rect -38 1398 -4 1432
rect 450 1398 484 1432
rect -38 904 -4 938
rect 450 904 484 938
rect -38 738 -4 772
rect 450 738 484 772
rect -38 244 -4 278
rect 450 244 484 278
<< locali >>
rect -170 1976 -110 2010
rect 576 1976 636 2010
rect -170 1945 -136 1976
rect 602 1945 636 1976
rect -40 1475 -6 1479
rect -54 1398 -38 1432
rect -4 1398 12 1432
rect 434 1398 450 1432
rect 484 1398 500 1432
rect -40 981 -6 984
rect 452 981 486 985
rect -54 904 -38 938
rect -4 904 12 938
rect 434 904 450 938
rect 484 904 500 938
rect -54 738 -38 772
rect -4 738 12 772
rect 434 738 450 772
rect 484 738 500 772
rect -40 691 -6 695
rect 452 692 486 695
rect -54 244 -38 278
rect -4 244 12 278
rect 434 244 450 278
rect 484 244 500 278
rect -40 197 -6 201
rect 452 198 486 201
rect -170 -269 -136 -243
rect 602 -269 636 -243
rect -170 -303 -110 -269
rect 576 -303 636 -269
<< viali >>
rect 195 2010 274 2014
rect 195 1976 274 2010
rect 195 1969 274 1976
rect -38 1398 -4 1432
rect 450 1398 484 1432
rect -38 904 -4 938
rect 450 904 484 938
rect -38 738 -4 772
rect 450 738 484 772
rect -38 244 -4 278
rect 450 244 484 278
<< metal1 >>
rect 183 2014 286 2020
rect 183 1969 195 2014
rect 274 1969 286 2014
rect 183 1963 286 1969
rect 436 1936 446 1938
rect 0 1935 43 1936
rect 396 1935 446 1936
rect 0 1884 446 1935
rect 0 1844 43 1884
rect 436 1880 446 1884
rect 502 1880 512 1938
rect -41 1485 -34 1668
rect 0 1485 42 1844
rect 108 1719 189 1766
rect 266 1721 342 1773
rect 360 1681 485 1683
rect 43 1485 83 1668
rect 180 1488 190 1669
rect 253 1488 263 1669
rect 360 1487 398 1681
rect 451 1674 485 1681
rect 451 1491 496 1674
rect 451 1487 489 1491
rect -34 1479 9 1485
rect 360 1482 489 1487
rect -50 1432 9 1479
rect -50 1398 -38 1432
rect -4 1398 9 1432
rect -50 1393 9 1398
rect -50 1392 0 1393
rect 107 1391 188 1438
rect 131 1346 159 1391
rect 254 1388 264 1440
rect 340 1388 350 1440
rect 451 1438 489 1482
rect 438 1432 496 1438
rect 438 1398 450 1432
rect 484 1398 496 1432
rect 438 1392 496 1398
rect 131 1318 316 1346
rect 86 1222 96 1274
rect 191 1222 201 1274
rect 288 1271 316 1318
rect 264 1224 345 1271
rect -42 1179 0 1181
rect -51 1178 0 1179
rect 43 1179 86 1181
rect 43 1178 87 1179
rect -60 984 -50 1178
rect 3 985 87 1178
rect 182 995 192 1176
rect 255 995 265 1176
rect 362 1174 496 1181
rect 357 998 440 1174
rect 492 998 496 1174
rect 357 991 491 998
rect 3 984 13 985
rect -50 938 8 984
rect -50 904 -38 938
rect -4 904 8 938
rect -50 894 8 904
rect 105 898 186 945
rect 451 944 489 985
rect 263 896 344 943
rect 438 938 496 944
rect 438 904 450 938
rect 484 904 496 938
rect 438 898 496 904
rect -52 772 8 784
rect -52 738 -38 772
rect -4 738 8 772
rect -52 697 8 738
rect 103 731 184 778
rect 257 732 346 783
rect 438 772 496 778
rect 438 738 450 772
rect 484 738 496 772
rect 438 732 496 738
rect -52 688 83 697
rect -62 506 -52 688
rect 2 506 83 688
rect -49 493 83 506
rect 180 503 190 684
rect 253 503 263 684
rect 446 682 493 732
rect 360 680 494 682
rect 360 504 440 680
rect 492 504 494 680
rect 360 499 494 504
rect 85 400 95 452
rect 190 400 200 452
rect 266 403 347 450
rect 287 361 322 403
rect 125 331 322 361
rect -49 278 8 291
rect 125 283 163 331
rect -49 244 -38 278
rect -4 244 8 278
rect -49 234 8 244
rect 108 236 189 283
rect 244 237 254 289
rect 349 237 359 289
rect 438 278 496 284
rect 438 244 450 278
rect 484 244 496 278
rect 438 238 496 244
rect -47 194 7 234
rect 446 198 496 238
rect -47 187 46 194
rect 386 187 396 198
rect -47 6 80 187
rect -47 -3 46 6
rect 179 4 189 185
rect 252 4 262 185
rect 357 4 396 187
rect 449 168 496 198
rect 449 4 491 168
rect 2 -208 46 -3
rect 108 -91 189 -44
rect 265 -91 346 -44
rect 424 -208 434 -206
rect 1 -279 434 -208
rect 351 -280 434 -279
rect 511 -280 521 -206
<< via1 >>
rect 446 1880 502 1938
rect 190 1488 253 1669
rect 398 1487 451 1681
rect 264 1388 340 1440
rect 96 1222 191 1274
rect -50 984 3 1178
rect 192 995 255 1176
rect 440 998 492 1174
rect -52 506 2 688
rect 190 503 253 684
rect 440 504 492 680
rect 95 400 190 452
rect 254 237 349 289
rect 189 4 252 185
rect 396 4 449 198
rect 434 -280 511 -206
<< metal2 >>
rect 446 1944 502 1948
rect 446 1938 503 1944
rect 502 1934 503 1938
rect 446 1878 447 1880
rect 446 1870 503 1878
rect 447 1868 503 1870
rect 405 1834 444 1837
rect -41 1795 444 1834
rect -41 1188 -2 1795
rect 405 1691 444 1795
rect 398 1681 451 1691
rect 190 1669 253 1679
rect 190 1478 253 1488
rect 398 1477 451 1487
rect 264 1440 340 1450
rect 264 1378 340 1388
rect 288 1346 316 1378
rect 131 1318 316 1346
rect 131 1284 159 1318
rect 96 1274 191 1284
rect 96 1214 191 1222
rect -50 1178 3 1188
rect 192 1176 255 1186
rect 192 985 255 995
rect 440 1175 498 1185
rect 440 987 498 997
rect -50 974 3 984
rect -41 698 -2 974
rect -52 688 2 698
rect -52 496 2 506
rect 190 684 253 694
rect -41 -121 -2 496
rect 190 493 253 503
rect 439 680 497 690
rect 439 492 497 502
rect 95 452 190 462
rect 95 390 190 400
rect 125 361 163 390
rect 125 331 322 361
rect 287 299 322 331
rect 254 289 349 299
rect 254 227 349 237
rect 396 198 449 208
rect 189 185 252 195
rect 189 -6 252 4
rect 396 -6 449 4
rect 405 -121 444 -6
rect -41 -160 444 -121
rect 434 -206 511 -196
rect 434 -290 511 -280
<< via2 >>
rect 447 1880 502 1934
rect 502 1880 503 1934
rect 447 1878 503 1880
rect 193 1489 251 1667
rect 193 997 251 1175
rect 440 1174 498 1175
rect 440 998 492 1174
rect 492 998 498 1174
rect 440 997 498 998
rect 193 503 251 681
rect 439 504 440 680
rect 440 504 492 680
rect 492 504 497 680
rect 439 502 497 504
rect 193 7 251 185
rect 445 -274 506 -213
<< metal3 >>
rect 446 1943 506 1944
rect 445 1939 506 1943
rect 437 1934 513 1939
rect 437 1878 447 1934
rect 503 1878 513 1934
rect 437 1873 513 1878
rect 191 1672 258 1679
rect 183 1667 261 1672
rect 183 1489 193 1667
rect 251 1489 261 1667
rect 183 1484 261 1489
rect 191 1180 258 1484
rect 445 1180 506 1873
rect 183 1175 261 1180
rect 183 997 193 1175
rect 251 997 261 1175
rect 183 992 261 997
rect 430 1175 508 1180
rect 430 997 440 1175
rect 498 997 508 1175
rect 430 992 508 997
rect 191 686 258 992
rect 183 681 261 686
rect 445 685 506 992
rect 183 503 193 681
rect 251 503 261 681
rect 183 498 261 503
rect 429 680 507 685
rect 429 502 439 680
rect 497 502 507 680
rect 191 190 258 498
rect 429 497 507 502
rect 183 185 261 190
rect 183 7 193 185
rect 251 7 261 185
rect 183 2 261 7
rect 445 -208 506 497
rect 435 -213 516 -208
rect 435 -274 445 -213
rect 506 -274 516 -213
rect 435 -279 516 -274
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1729246168
transform 1 0 21 0 1 97
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1729246168
transform 1 0 425 0 1 1579
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1729246168
transform 1 0 425 0 1 1085
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_3
timestamp 1729246168
transform 1 0 425 0 1 591
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_4
timestamp 1729246168
transform 1 0 425 0 1 97
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_5
timestamp 1729246168
transform 1 0 21 0 1 1579
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_6
timestamp 1729246168
transform 1 0 21 0 1 1085
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_7
timestamp 1729246168
transform 1 0 21 0 1 591
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_VQXX5L  sky130_fd_pr__pfet_01v8_VQXX5L_0
timestamp 1729273948
transform 1 0 223 0 1 591
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_VQXX5L  sky130_fd_pr__pfet_01v8_VQXX5L_1
timestamp 1729273948
transform 1 0 223 0 1 97
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_VQXX5L  sky130_fd_pr__pfet_01v8_VQXX5L_2
timestamp 1729273948
transform 1 0 223 0 1 1085
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_VQXX5L  sky130_fd_pr__pfet_01v8_VQXX5L_3
timestamp 1729273948
transform 1 0 223 0 1 1579
box -223 -200 223 200
<< labels >>
flabel metal3 217 836 217 836 0 FreeSans 480 0 0 0 D5
port 0 nsew
flabel metal1 144 1364 144 1364 0 FreeSans 480 0 0 0 VIP
port 1 nsew
flabel metal2 299 1364 299 1364 0 FreeSans 480 0 0 0 VIN
port 2 nsew
flabel metal2 136 1819 136 1819 0 FreeSans 480 0 0 0 D6
port 3 nsew
flabel metal3 480 1780 480 1780 0 FreeSans 480 0 0 0 OUT
port 4 nsew
flabel viali 229 1989 229 1989 0 FreeSans 480 0 0 0 VDD
port 5 nsew
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1729397805
<< viali >>
rect -2179 3129 -2137 3163
<< metal1 >>
rect -1631 4011 -1180 4062
rect -1231 3407 -1180 4011
rect -1648 3211 -1638 3266
rect -1583 3211 -1573 3266
rect -2191 3163 -2124 3175
rect -2191 3129 -2179 3163
rect -2137 3129 -2124 3163
rect -2191 3121 -2124 3129
rect -2178 2971 -2137 3121
rect -1602 2820 -297 2821
rect -1602 2819 -294 2820
rect -1602 2785 -249 2819
rect -371 2734 -249 2785
rect -371 2698 -247 2734
rect -371 2696 -325 2698
rect -371 2676 -286 2696
rect -283 2676 -247 2698
rect -371 2641 -247 2676
rect -371 2640 -266 2641
rect -1658 1820 -1600 1865
rect -552 1820 -494 2032
rect -1658 1762 -494 1820
<< via1 >>
rect -1638 3211 -1583 3266
<< metal2 >>
rect -1638 3266 -1583 3276
rect -1650 3223 -1638 3262
rect -1130 3262 -1091 3285
rect -1583 3223 -1090 3262
rect -1130 3212 -1091 3223
rect -1638 3201 -1583 3211
<< metal3 >>
rect -646 2675 -586 3289
rect -1804 2408 -1748 2555
rect -1816 2348 -1748 2408
rect -1815 2347 -1748 2348
rect -1804 2346 -1748 2347
use nmos89  nmos89_0 ~/opamp/mag/nmos89
timestamp 1729231471
transform 1 0 -2602 0 -1 4005
box -177 -131 1107 884
use nmoscs  nmoscs_0 ~/opamp/mag/nmoscs
timestamp 1729266392
transform 1 0 -2446 0 1 2400
box -409 -811 1089 721
use pmos67  pmos67_0 ~/opamp/mag/pmos67
timestamp 1729350307
transform 0 -1 704 1 0 3040
box -206 -342 672 2046
use pmoscs  pmoscs_0 ~/opamp/mag/pmoscs
timestamp 1729348601
transform 0 -1 734 1 0 2034
box -238 -820 833 2087
<< labels >>
flabel metal1 -2158 3068 -2158 3068 0 FreeSans 800 0 0 0 GND
port 0 nsew
flabel metal2 -1448 3242 -1448 3242 0 FreeSans 800 0 0 0 D8
port 1 nsew
flabel metal1 -1212 4032 -1212 4032 0 FreeSans 800 0 0 0 OUT
port 2 nsew
flabel metal3 -620 2850 -620 2850 0 FreeSans 800 0 0 0 D5
port 3 nsew
flabel metal1 -324 2756 -324 2756 0 FreeSans 800 0 0 0 D2
port 4 nsew
flabel metal1 -960 1798 -960 1798 0 FreeSans 800 0 0 0 D1
port 5 nsew
<< end >>

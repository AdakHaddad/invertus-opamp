magic
tech sky130A
magscale 1 2
timestamp 1729180798
<< pwell >>
rect -425 -410 425 410
<< nmos >>
rect -229 -200 -29 200
rect 29 -200 229 200
<< ndiff >>
rect -287 188 -229 200
rect -287 -188 -275 188
rect -241 -188 -229 188
rect -287 -200 -229 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 229 188 287 200
rect 229 -188 241 188
rect 275 -188 287 188
rect 229 -200 287 -188
<< ndiffc >>
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
<< psubdiff >>
rect -389 340 -293 374
rect 293 340 389 374
rect -389 278 -355 340
rect 355 278 389 340
rect -389 -340 -355 -278
rect 355 -340 389 -278
rect -389 -374 -293 -340
rect 293 -374 389 -340
<< psubdiffcont >>
rect -293 340 293 374
rect -389 -278 -355 278
rect 355 -278 389 278
rect -293 -374 293 -340
<< poly >>
rect -229 272 -29 288
rect -229 238 -213 272
rect -45 238 -29 272
rect -229 200 -29 238
rect 29 272 229 288
rect 29 238 45 272
rect 213 238 229 272
rect 29 200 229 238
rect -229 -238 -29 -200
rect -229 -272 -213 -238
rect -45 -272 -29 -238
rect -229 -288 -29 -272
rect 29 -238 229 -200
rect 29 -272 45 -238
rect 213 -272 229 -238
rect 29 -288 229 -272
<< polycont >>
rect -213 238 -45 272
rect 45 238 213 272
rect -213 -272 -45 -238
rect 45 -272 213 -238
<< locali >>
rect -389 340 -293 374
rect 293 340 389 374
rect -389 278 -355 340
rect 355 278 389 340
rect -229 238 -213 272
rect -45 238 -29 272
rect 29 238 45 272
rect 213 238 229 272
rect -275 188 -241 204
rect -275 -204 -241 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 241 188 275 204
rect 241 -204 275 -188
rect -229 -272 -213 -238
rect -45 -272 -29 -238
rect 29 -272 45 -238
rect 213 -272 229 -238
rect -389 -340 -355 -278
rect 355 -340 389 -278
rect -389 -374 -293 -340
rect 293 -374 389 -340
<< viali >>
rect -213 238 -45 272
rect 45 238 213 272
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect -213 -272 -45 -238
rect 45 -272 213 -238
<< metal1 >>
rect -225 272 -33 278
rect -225 238 -213 272
rect -45 238 -33 272
rect -225 232 -33 238
rect 33 272 225 278
rect 33 238 45 272
rect 213 238 225 272
rect 33 232 225 238
rect -281 188 -235 200
rect -281 -188 -275 188
rect -241 -188 -235 188
rect -281 -200 -235 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 235 188 281 200
rect 235 -188 241 188
rect 275 -188 281 188
rect 235 -200 281 -188
rect -225 -238 -33 -232
rect -225 -272 -213 -238
rect -45 -272 -33 -238
rect -225 -278 -33 -272
rect 33 -238 225 -232
rect 33 -272 45 -238
rect 213 -272 225 -238
rect 33 -278 225 -272
<< properties >>
string FIXED_BBOX -372 -357 372 357
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 1 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

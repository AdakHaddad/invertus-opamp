magic
tech sky130A
timestamp 1729264637
<< nmos >>
rect -50 -21 50 21
<< ndiff >>
rect -79 15 -50 21
rect -79 -15 -73 15
rect -56 -15 -50 15
rect -79 -21 -50 -15
rect 50 15 79 21
rect 50 -15 56 15
rect 73 -15 79 15
rect 50 -21 79 -15
<< ndiffc >>
rect -73 -15 -56 15
rect 56 -15 73 15
<< poly >>
rect -50 57 50 65
rect -50 40 -42 57
rect 42 40 50 57
rect -50 21 50 40
rect -50 -40 50 -21
rect -50 -57 -42 -40
rect 42 -57 50 -40
rect -50 -65 50 -57
<< polycont >>
rect -42 40 42 57
rect -42 -57 42 -40
<< locali >>
rect -50 40 -42 57
rect 42 40 50 57
rect -73 15 -56 23
rect -73 -23 -56 -15
rect 56 15 73 23
rect 56 -23 73 -15
rect -50 -57 -42 -40
rect 42 -57 50 -40
<< viali >>
rect -42 40 42 57
rect -73 -15 -56 15
rect 56 -15 73 15
rect -42 -57 42 -40
<< metal1 >>
rect -48 57 48 60
rect -48 40 -42 57
rect 42 40 48 57
rect -48 37 48 40
rect -76 15 -53 21
rect -76 -15 -73 15
rect -56 -15 -53 15
rect -76 -21 -53 -15
rect 53 15 76 21
rect 53 -15 56 15
rect 73 -15 76 15
rect 53 -21 76 -15
rect -48 -40 48 -37
rect -48 -57 -42 -40
rect 42 -57 48 -40
rect -48 -60 48 -57
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.420 l 1 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
